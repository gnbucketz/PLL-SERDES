`timescale 1ns / 1ps

module Frequency_Divider#(
parameter n = 1
//1 d FF = divide 2, 2 d FF = divide 4, 3 d FF = divide by 8
)(
input clk, input rst, input d1, input d2, input d3, input qn1, input qn2, input qn3, output reg q1, output reg q2, output reg q3

   
   
    );
endmodule
